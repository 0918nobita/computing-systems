module OR(a, b, OUT);
    input a;
    input b;
    output OUT;

    assign OUT = a | b;
endmodule
