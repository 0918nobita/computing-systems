module main ();
    initial $display("Hello, world!");
endmodule
